module switch_sva(
);

endmodule
