bind switch switch_sva sva_inst(
*.
);

endmodule
